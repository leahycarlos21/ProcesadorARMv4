module restador# (parameter size = 32)(input logic [size-1:0] a, b,
											output logic [size-1:0] result);
											

																			
assign result = a-b;




endmodule 