module xor_# (parameter size = 4)(input logic [size-1:0] a, b,
				output logic [size-1:0] c);
assign c = a ^ b;
endmodule